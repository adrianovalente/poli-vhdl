library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

entity calc is
  port(
    time_in: in integer range 0 to 24000;
    alg0, alg1, alg2, color: out std_logic_vector(3 downto 0)
  );
end calc;

architecture seila of calc is
  signal dist: integer range 0 to 512;
  signal first, second: integer range 0 to 512;
begin
  if time_in<20 then
    color <= "1111";
  else
    if time_in<40 then
      color <= "1011";
    else
      color <= "1010";
    end if;
  end if;
  dist <= time_in/58;
  alg0 <= std_logic_vector(to_unsigned(dist mod 10, alg0'length));
  first <= dist/10;
  alg1 <= std_logic_vector(to_unsigned(first mod 10, alg1'length));
  second <= first/10;
  alg2 <= std_logic_vector(to_unsigned(second mod 10, alg2'length));
end seila;
